`ifndef GUARD_UART_DEFINE__SV
`define GUARD_UART_DEFINE__SV
     
     `ifndef UART_DATA_WIDTH
          `define UART_DATA_WIDTH 14
     `endif
`endif
